magic
tech scmos
timestamp 1445617567
<< pwell >>
rect -5 -2 11 10
<< nwell >>
rect -3 20 9 32
<< polysilicon >>
rect 2 24 4 26
rect 2 9 4 21
rect 2 4 4 6
<< ndiffusion >>
rect 1 6 2 9
rect 4 6 5 9
<< pdiffusion >>
rect 1 21 2 24
rect 4 21 5 24
<< metal1 >>
rect 1 28 9 32
rect -3 24 1 28
rect 5 17 9 20
rect -7 13 -2 17
rect 5 13 15 17
rect 5 10 9 13
rect -3 2 1 6
rect 1 -2 9 2
<< ntransistor >>
rect 2 6 4 9
<< ptransistor >>
rect 2 21 4 24
<< polycontact >>
rect -2 13 2 17
<< ndcontact >>
rect -3 6 1 10
rect 5 6 9 10
<< pdcontact >>
rect -3 20 1 24
rect 5 20 9 24
<< psubstratepcontact >>
rect -3 -2 1 2
<< nsubstratencontact >>
rect -3 28 1 32
<< labels >>
rlabel metal1 -5 15 -5 15 3 IN
rlabel metal1 9 15 9 15 7 OUT
rlabel metal1 3 30 3 30 5 VDD
rlabel metal1 3 0 3 0 1 GND
<< end >>
